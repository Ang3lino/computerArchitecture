LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY MEMORIA_PROGRAMA IS
	-- VALORES GENERICOS DE LA MEMORIA DE PROGRAMA DEL ESCOMIPS
	GENERIC(
		BITS_A : INTEGER := 25;
		BITS_D : INTEGER := 16);

	-- PUERTOS DE ENTRADA (BUS DE DIRECCIONES 'A')
	-- Y SALIDA (BUS DE DIRECCIONES 'D')
    PORT ( A : IN STD_LOGIC_VECTOR (BITS_D - 1 DOWNTO 0);
           D : OUT STD_LOGIC_VECTOR (BITS_A - 1 DOWNTO 0));
END MEMORIA_PROGRAMA;

ARCHITECTURE FUNCIONAMIENTO OF MEMORIA_PROGRAMA IS
	-- C�DIGOS DE OPERACI�N DE CADA UNA DE LAS INSTRUCCIONES.
	CONSTANT OPCODE_TIPOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000"; -- OPERACIONES _00 (TIPO R)
	CONSTANT OPCODE_LI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
	CONSTANT OPCODE_LWI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
	CONSTANT OPCODE_SWI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
	CONSTANT OPCODE_SW		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
	CONSTANT OPCODE_ADDI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
	CONSTANT OPCODE_SUBI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
	CONSTANT OPCODE_ANDI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
	CONSTANT OPCODE_ORI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
	CONSTANT OPCODE_XORI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
	CONSTANT OPCODE_NANDI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
	CONSTANT OPCODE_NORI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
	CONSTANT OPCODE_XNORI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
	CONSTANT OPCODE_BEQI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
	CONSTANT OPCODE_BNEI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
	CONSTANT OPCODE_BLTI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
	CONSTANT OPCODE_BLETI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
	CONSTANT OPCODE_BGTI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
	CONSTANT OPCODE_BGETI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
	CONSTANT OPCODE_B		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
	CONSTANT OPCODE_CALL	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10100";
	CONSTANT OPCODE_RET		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10101";
	CONSTANT OPCODE_NOP		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10110";
	CONSTANT OPCODE_LW 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
	-- ...

	-- C�DIGOS DE VARIACI�N DE LA OPERACI�N ADD
	CONSTANT FUNCODE_ADD	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	CONSTANT FUNCODE_SUB	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";

	-- REGISTROS	
	CONSTANT R_00	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	CONSTANT R_01	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
	CONSTANT R_02	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
	CONSTANT R_03	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
	CONSTANT R_04	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
	CONSTANT R_05	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";
	CONSTANT R_06	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
	CONSTANT R_07	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
	CONSTANT R_08	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
	CONSTANT R_09	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
	CONSTANT R_10	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
	CONSTANT R_11	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";
	CONSTANT R_12	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";
	CONSTANT R_13	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101";
	CONSTANT R_14	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1110";
	CONSTANT R_15	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111";

	-- SIN USAR	
	CONSTANT SIN_USO		: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	
	-- DEFIINICI�N DEL TIPO DE DATO MEMORIA
	TYPE MEMORIA IS ARRAY (0 TO 2 ** BITS_A - 1) 
		OF STD_LOGIC_VECTOR(BITS_A - 1 DOWNTO 0); 

	-- DECLARACI�N DE UNA MEMORIA ROM CON EL PROGRAMA DE EJEMPLO.
	CONSTANT ROM : MEMORIA := (
		OPCODE_LI 	 & R_00 	& X"0001",
		OPCODE_LI 	 & R_01 	& X"0007",
		OPCODE_TIPOR & R_01 	& R_01 & R_00 & SIN_USO & FUNCODE_ADD,
		OPCODE_SWI 	 & R_01 	& X"0005",
		OPCODE_B 	 & SIN_USO 	& X"0002",
		OTHERS => (OTHERS => '0'));

BEGIN

	-- LECTURA ASINCRONA DE LA MEMORIA.
	D <= ROM(CONV_INTEGER(A));

END FUNCIONAMIENTO;

