----------------------------------------------------------------------------------
-- Authors:
		-- Lpez Manriquez ngel
		-- Maya Rocha Luis Emmanuel
		-- Vazquez Moreno Marcos Oswaldo
-- Create Date:    17:22:07 10/06/2018 
-- Module Name:    Memory - Behavioral 
-- Project Name: ProgramMem
--
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;


entity program_memory is
	Generic (BADDR: Integer:=16;
			  BDATA: Integer:=25 );
    Port ( A : in  STD_LOGIC_VECTOR (BADDR-1 downto 0);
		   D : out  STD_LOGIC_VECTOR (BDATA-1 downto 0)
	);
end program_memory;

architecture BEHAVIOR of program_memory is
-- Operation codes
	CONSTANT OPCODE_TIPOR 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
	CONSTANT OPCODE_LI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
	CONSTANT OPCODE_LWI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
	CONSTANT OPCODE_SWI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
	CONSTANT OPCODE_SW   	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
	CONSTANT OPCODE_ADDI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
	CONSTANT OPCODE_SUBI		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
	CONSTANT OPCODE_ANDI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
	CONSTANT OPCODE_ORI 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
	CONSTANT OPCODE_XORI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
	CONSTANT OPCODE_NANDI	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
	CONSTANT OPCODE_NORI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
	CONSTANT OPCODE_XNORI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
	CONSTANT OPCODE_BEQI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
	CONSTANT OPCODE_BNEI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
	CONSTANT OPCODE_BLTI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
	CONSTANT OPCODE_BLETI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";
	CONSTANT OPCODE_BGTI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10001";
	CONSTANT OPCODE_BGETI 	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10010";
	CONSTANT OPCODE_B   	   : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10011";
	CONSTANT OPCODE_CALL		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10100";
	CONSTANT OPCODE_RET		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10101";
	CONSTANT OPCODE_NOP  	: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10110";
	CONSTANT OPCODE_LW 		: STD_LOGIC_VECTOR(4 DOWNTO 0) := "10111";

-- R Instructions' functions
	CONSTANT FUN_ADD			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	CONSTANT FUN_SUB			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";	
	CONSTANT FUN_AND			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
	CONSTANT FUN_OR			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";	
	CONSTANT FUN_XOR			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
	CONSTANT FUN_NAND	  	   : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";	
	CONSTANT FUN_NOR			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
	CONSTANT FUN_XNOR	   	: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";	
	CONSTANT FUN_NOT			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
	CONSTANT FUN_SLL			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";	
	CONSTANT FUN_SRL			: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";	

--Process registers:
	CONSTANT R0					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
	CONSTANT R1					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
	CONSTANT R2					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
	CONSTANT R3					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
	CONSTANT R4					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
	CONSTANT R5					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";	
	CONSTANT R6					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0110";
	CONSTANT R7					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0111";
	CONSTANT R8					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1000";
	CONSTANT R9					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1001";
	CONSTANT R10				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1010";
	CONSTANT R11				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1011";	
	CONSTANT R12				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1100";
	CONSTANT R13				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1101";	
	CONSTANT R14				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1110";
	CONSTANT R15				: STD_LOGIC_VECTOR(3 DOWNTO 0) := "1111";	
	CONSTANT SU					: STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";

	TYPE ARR IS ARRAY (0 TO 2**BADDR - 1) OF STD_LOGIC_VECTOR(D'RANGE); 
	CONSTANT ROM : ARR := (
	--Instructions:
		OPCODE_LI&R0&X"0001",
		OPCODE_LI&R1&X"0007",
		OPCODE_TIPOR&R1&R1&R0&SU&FUN_ADD,
		OPCODE_SWI&R1&X"0005",
		OPCODE_B&SU&X"0002",
		OTHERS=>(OTHERS=>'0')
	);

begin

	D <= ROM( CONV_INTEGER(A) );
end BEHAVIOR;