
library IEEE;
LIBRARY WORK;

use IEEE.STD_LOGIC_1164.ALL;
USE WORK.components.ALL;

ENTITY main IS
	PORT ( 
		CLK	: IN STD_LOGIC;
		CLR	: IN STD_LOGIC;
		datain: inout std_logic_vector(15 downto 0)
	);
END main;

ARCHITECTURE ESCOMIPS OF main IS

	signal clk_reduced : STD_LOGIC;
    signal SAL_ALU : STD_LOGIC_VECTOR(15 DOWNTO 0);
	signal wd: std_logic;
	signal BANDAS : STD_LOGIC_VECTOR(3 DOWNTO 0);


    --SIGNAL CLK 	:	STD_LOGIC;
    SIGNAL SALIDA_CONTROL : STD_LOGIC_VECTOR(19 DOWNTO 0);
    SIGNAL SALIDA_PILA : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_SOP1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_SOP2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_SDMP : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_MEM_PROG : STD_LOGIC_VECTOR(24 DOWNTO 0);
    SIGNAL READ_DATA1 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL READ_DATA2 : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL READ_REGISTER2 : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL WRITE_DATA : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_SR : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_SEXT : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL BANDERAS : STD_LOGIC_VECTOR(3 DOWNTO 0);
    SIGNAL SALIDA_ALU : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_SDMD : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_RAM : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_EXT_DIR : STD_LOGIC_VECTOR(15 DOWNTO 0);
    SIGNAL SALIDA_EXT_SIG : STD_LOGIC_VECTOR(15 DOWNTO 0);

    constant logic_one: std_logic := '1';

BEGIN

	datain <= read_data2;

	DIV : DIVISOR PORT MAP(
		OSC_CLK		=> 	CLK,
		CLR			=>	CLR,
		CLK			=>	clk_reduced
	);

	SAL_ALU <= SALIDA_ALU;
	WD		<= SALIDA_CONTROL(1);
	BANDAS <= SALIDA_CONTROL(6 DOWNTO 3);

	MEM_PROG : program_memory PORT MAP(
		A => SALIDA_PILA,
        D => SALIDA_MEM_PROG,
        clk => clk
	);
	
	SALIDA_SOP1 <= SALIDA_PILA WHEN (SALIDA_CONTROL(8) = '1') ELSE READ_DATA1;
	
	SALIDA_SDMP <= SALIDA_SR WHEN (SALIDA_CONTROL(16) = '1') ELSE SALIDA_MEM_PROG(15 DOWNTO 0);

	PILA_HW	: stack PORT MAP(
		CLK 	=> CLK_reduced,
		CLR 	=> CLR,
		WPC	=> SALIDA_CONTROL(17),
		UP		=> SALIDA_CONTROL(19),
		DW		=> SALIDA_CONTROL(18),
		D 		=> SALIDA_SDMP,
		Q		=> SALIDA_PILA
	); --

	READ_REGISTER2 <= SALIDA_MEM_PROG(19 DOWNTO 16) WHEN (SALIDA_CONTROL(15) = '1') ELSE 
							SALIDA_MEM_PROG(11 DOWNTO 8);

	WRITE_DATA <= SALIDA_SR WHEN (SALIDA_CONTROL(14) = '1') ELSE 
						SALIDA_MEM_PROG(15 DOWNTO 0);
	
	ARCH_REG : file_register PORT MAP(
		READ_REGISTER_1 => SALIDA_MEM_PROG(15 DOWNTO 12),
		READ_REGISTER_2 => READ_REGISTER2,
		WRITE_REGISTER => SALIDA_MEM_PROG(19 DOWNTO 16),
		SHAMT				=> SALIDA_MEM_PROG(7 DOWNTO 4),
		WRITE_DATA 		=> WRITE_DATA,
		CLK				=> CLK_reduced,
		SHE 				=> SALIDA_CONTROL(13),
		DIR				=> SALIDA_CONTROL(12),
		We					=> SALIDA_CONTROL(11),
		READ_DATA_1		=> READ_DATA1,
		READ_DATA_2		=> READ_DATA2
	); --


	SALIDA_EXT_DIR <= X"0"&SALIDA_MEM_PROG(11 DOWNTO 0);
	SALIDA_EXT_SIG <= X"F"&SALIDA_MEM_PROG(11 DOWNTO 0) WHEN (SALIDA_MEM_PROG(11) = '1')
							ELSE X"0"&SALIDA_MEM_PROG(11 DOWNTO 0);

	SALIDA_SEXT <= SALIDA_EXT_DIR WHEN (SALIDA_CONTROL(9) = '1') ELSE
						SALIDA_EXT_SIG;


	SALIDA_SOP2 <= SALIDA_SEXT WHEN (SALIDA_CONTROL(7) = '1') ELSE 
                        READ_DATA2;
    
	MEM_DATOS : memoria_datos PORT MAP(
		WD		=> SALIDA_CONTROL(1),
		CLK	    => CLK_reduced,
		ADR 	=> SALIDA_SDMD,
		bus_datos_entrada	=> READ_DATA2,
        bus_datos_salida 	=> SALIDA_RAM,
        rd => logic_one
	); --

	ALU_MIPS : ALU PORT MAP(
		A 	=> SALIDA_SOP1,
		B 	=> SALIDA_SOP2,
		ALUOP	=> SALIDA_CONTROL(6 DOWNTO 3),
		flags => BANDERAS,
		ans => SALIDA_ALU
	); -- 

	SALIDA_SDMD <= SALIDA_MEM_PROG(15 DOWNTO 0) WHEN (SALIDA_CONTROL(2) = '1') ELSE
						SALIDA_ALU;

	SALIDA_SR <= SALIDA_ALU WHEN (SALIDA_CONTROL(1) = '1') ELSE
					SALIDA_RAM;

	UNIDAD_CTRL : CONTROL PORT MAP(
		OPCODE 	=>	SALIDA_MEM_PROG(24 DOWNTO 20),
		FUNCODE	=>	SALIDA_MEM_PROG(3 DOWNTO 0),
		flags	=>	BANDERAS,
		CLK		=>	CLK_reduced,
		CLR		=>	CLR,
		LF		=>	SALIDA_CONTROL(10),
		s 	=>	SALIDA_CONTROL
	); --

END ESCOMIPS;

